module tb_adder();

	reg clk = 0;
	reg scan_clk = 0;
	reg reset = 0;
	reg clb_scan_in, clb_scan_en, conn_scan_in, conn_scan_en;

	reg start_fpga_clk = 0;	wire clb_scan_out, conn_scan_out;
	wire [19:0] fpga_io;
    reg [19:0] is_fpga_input = {4'b0111, 4'b1101, 4'b0111, 4'b0001, 4'b1110};

    reg [19:0] fpga_input=20'h0;

	reg [5:0] a = 5'b00011;
	reg [5:0] b = 5'b00011;
    
    genvar i;
	generate
		for(i = 0; i < 20; i = i + 1) begin
			assign fpga_io[i] = is_fpga_input[i] ? fpga_input[i] : 1'bz;
		end
	endgenerate
    
    //assign fpga_io[14] = tristate ? fpga_reset_in : 1'bz;
    
    chip inst_chip(
		.clk(clk),
		.scan_clk(scan_clk),
		.fpga_io(fpga_io),
		.clb_scan_in(clb_scan_in),
		.clb_scan_out(clb_scan_out),
		.clb_scan_en(clb_scan_en),
		.conn_scan_in(conn_scan_in),
		.conn_scan_out(conn_scan_out),
		.conn_scan_en(conn_scan_en),
		.reset(reset)
	);

	initial begin
		clk = 0; scan_clk = 0; reset = 0; clb_scan_in = 0; clb_scan_en = 0; conn_scan_in = 0; conn_scan_en = 0;
	end

	always begin
		#5 scan_clk = ~scan_clk;
	end
    always @(*) begin
		if (start_fpga_clk)
			clk = scan_clk;
		else
			clk = 0;
	end	
    initial begin
		$dumpfile("tb_adder.vcd");
		$dumpvars(0, tb_adder);
    		#10 clb_scan_en <= 1; clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_en <= 0;
		#10 conn_scan_en <= 1; conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_en <= 0; start_fpga_clk <= 1;
		#10 reset <= 1;
		#10 reset <= 0;
		// out[0] = sum[3] in[1]=b[4] in[3]=b[3] in[4]=a[3] out[5]=sum[4] out[6]=sum[5] out[7]=sum[6]
 		// in[8] = b[5] in[9]=a[4] in[10]=a[2] out[11]=sum[0] in[12]=a[5] out[13]=sum[1] in[14]=a[0]
 		// in[15] = b[1] in[16]=a[1] in[17]=b[0] in[18]=b[2] out[19]=sum[2]
 		

 		// sum = 6'b000100
 		
 		#10 fpga_input[14] <= a[0]; fpga_input[16] <= a[1]; fpga_input[10] <= a[2]; fpga_input[4] <= a[3]; fpga_input[12] <= a[5]; 
 		fpga_input[17] <= b[0]; fpga_input[15] <= b[1]; fpga_input[18] <= b[2]; fpga_input[3] <= b[3]; fpga_input[8] <= b[5]; 
 
		#5000 $finish;
	 end
endmodule