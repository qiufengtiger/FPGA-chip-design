module tb_blink();
	reg clk = 0;
	reg scan_clk = 0;
	reg reset = 0;
	reg clb_scan_in, clb_scan_en, conn_scan_in, conn_scan_en;

	reg start_fpga_clk = 0;	wire clb_scan_out, conn_scan_out;
	reg [19:0] fpga_in = 0;
	wire [19:0] fpga_out;

	fpga_core inst_test_fpga_core(
		.clk(clk),
		.scan_clk(scan_clk),
		.fpga_in(fpga_in),
		.fpga_out(fpga_out),
		.clb_scan_in(clb_scan_in),
		.clb_scan_out(clb_scan_out),
		.clb_scan_en(clb_scan_en),
		.conn_scan_in(conn_scan_in),
		.conn_scan_out(conn_scan_out),
		.conn_scan_en(conn_scan_en),
		.reset(reset)
	);

	initial begin
		clk = 0; scan_clk = 0; reset = 0; clb_scan_in = 0; clb_scan_en = 0; conn_scan_in = 0; conn_scan_en = 0;
	end

	always begin
    #10
        if (~start_fpga_clk)
            scan_clk = ~scan_clk;
        else
            scan_clk = 0;
    end
	always begin
    #10
		if (start_fpga_clk)
			clk = ~clk;
		else
			clk = 0;
	end
	initial begin
		$dumpfile("tb_blink.vcd");
		$dumpvars(0, tb_blink);
		#10 clb_scan_en <= 1; clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b0;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_in <= 1'b1;
		#20 clb_scan_en <= 0;
		#20 conn_scan_en <= 1; conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b1;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_in <= 1'b0;
		#20 conn_scan_en <= 0; start_fpga_clk <= 1;
		#20 reset <= 1;
		#20 reset <= 0;
		#10 fpga_in[14] = 1'b1;
 		#10 fpga_in[14] = 1'b0;
 
		#100680 $finish;
	 end
endmodule