module blink_tb();
	reg clk = 0;
	reg scan_clk = 0;
	reg reset = 0;
	reg clb_scan_in, clb_scan_en, conn_scan_in, conn_scan_en;

	wire clb_scan_out, conn_scan_out;
	wire [19:0] fpga_in, fpga_out;

	fpga_core inst_test_fpga_core(
		.clk(clk),
		.scan_clk(scan_clk),
		.fpga_in(fpga_in),
		.fpga_out(fpga_out),
		.clb_scan_in(clb_scan_in),
		.clb_scan_out(clb_scan_out),
		.clb_scan_en(clb_scan_en),
		.conn_scan_in(conn_scan_in),
		.conn_scan_out(conn_scan_out),
		.conn_scan_en(conn_scan_en),
		.reset(reset)
	);

	initial begin
		clk = 0; scan_clk = 0; reset = 0; clb_scan_in = 0; clb_scan_en = 0; conn_scan_in = 0; conn_scan_en = 0;
	end

	always begin
		#5 scan_clk = ~scan_clk;
	end
	initial begin
		$dumpfile("blink_tb.vcd");
		$dumpvars(0, blink_tb);
		$dumpon;

		#10 clb_scan_en <= 1; clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b1;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_in <= 1'b0;
		#10 clb_scan_en <= 0
		#10 conn_scan_en <= 1; conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b1;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_in <= 1'b0;
		#10 conn_scan_en <= 0
		#10 fpga_in[14] = 1'b1; 
		#50440 $finish;
	 end
endmodule